<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-17.1889,17.8889,61.3889,-64.0667</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-3.5,-24.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>31.5,-24</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>6 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>BE_JKFF_LOW_NT</type>
<position>18.5,-24</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>3 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>BE_JKFF_LOW_NT</type>
<position>6,-24</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>4 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-3.5,-16.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>49,-30</position>
<input>
<ID>N_in3</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>11,-29</position>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>24.5,-29</position>
<input>
<ID>N_in3</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>BE_JKFF_LOW_NT</type>
<position>44.5,-24</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>38.5,-29</position>
<input>
<ID>N_in3</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>21.5,-6</position>
<gparam>LABEL_TEXT 4-Bit Asynchronous Counter</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-24.5,0.5,-24</points>
<intersection>-24.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-24,3,-24</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-24.5,0.5,-24.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-16.5,40,-16.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>1.5 5</intersection>
<intersection>13.5 10</intersection>
<intersection>26.5 9</intersection>
<intersection>40 17</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1.5,-26,1.5,-16.5</points>
<intersection>-26 7</intersection>
<intersection>-22 15</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>1.5,-26,3,-26</points>
<connection>
<GID>4</GID>
<name>K</name></connection>
<intersection>1.5 5</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>26.5,-26,26.5,-16.5</points>
<intersection>-26 19</intersection>
<intersection>-22 13</intersection>
<intersection>-16.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>13.5,-26,13.5,-16.5</points>
<intersection>-26 11</intersection>
<intersection>-22 14</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>13.5,-26,15.5,-26</points>
<connection>
<GID>3</GID>
<name>K</name></connection>
<intersection>13.5 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>26.5,-22,28.5,-22</points>
<connection>
<GID>2</GID>
<name>J</name></connection>
<intersection>26.5 9</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>13.5,-22,15.5,-22</points>
<connection>
<GID>3</GID>
<name>J</name></connection>
<intersection>13.5 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>1.5,-22,3,-22</points>
<connection>
<GID>4</GID>
<name>J</name></connection>
<intersection>1.5 5</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>40,-26,40,-16.5</points>
<intersection>-26 20</intersection>
<intersection>-22 21</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>26.5,-26,28.5,-26</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>26.5 9</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>40,-26,41.5,-26</points>
<connection>
<GID>9</GID>
<name>K</name></connection>
<intersection>40 17</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>40,-22,41.5,-22</points>
<connection>
<GID>9</GID>
<name>J</name></connection>
<intersection>40 17</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-28,24.5,-22</points>
<connection>
<GID>8</GID>
<name>N_in3</name></connection>
<intersection>-24 2</intersection>
<intersection>-22 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-24,28.5,-24</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-22,24.5,-22</points>
<connection>
<GID>3</GID>
<name>Q</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-28,11,-22</points>
<connection>
<GID>7</GID>
<name>N_in3</name></connection>
<intersection>-24 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,-24,15.5,-24</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>9,-22,11,-22</points>
<connection>
<GID>4</GID>
<name>Q</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-29,49,-22</points>
<connection>
<GID>6</GID>
<name>N_in3</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-22,49,-22</points>
<connection>
<GID>9</GID>
<name>Q</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-28,38.5,-22</points>
<connection>
<GID>10</GID>
<name>N_in3</name></connection>
<intersection>-24 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-24,41.5,-24</points>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34.5,-22,38.5,-22</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>