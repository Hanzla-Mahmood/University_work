<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.93846,12.3255,83.5383,-72.7819</PageViewport>
<gate>
<ID>2</ID>
<type>AE_OR4</type>
<position>88.5,-27</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>12 </input>
<input>
<ID>IN_3</ID>13 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>94,-27</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>62.5,-10.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND3</type>
<position>62.5,-22.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>62.5,-33.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND3</type>
<position>62.5,-45.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>13.5,-6.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>14,-11</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>13.5,-18.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>13.5,-28</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>13,-36</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>12.5,-47</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>28.5,-7.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>27,-11.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>8.5,-6</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>8,-11</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>7,-18.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>8,-27</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>7.5,-35.5</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>6.5,-46</position>
<gparam>LABEL_TEXT I4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92.5,-27,93,-27</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>4</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-7.5,21,-6.5</points>
<intersection>-7.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-7.5,26.5,-7.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection>
<intersection>24 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-6.5,21,-6.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-31.5,24,-7.5</points>
<intersection>-31.5 4</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-31.5,59.5,-31.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection>
<intersection>36.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>36.5,-43.5,36.5,-31.5</points>
<intersection>-43.5 6</intersection>
<intersection>-31.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>36.5,-43.5,59.5,-43.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>36.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-11.5,21,-11</points>
<intersection>-11.5 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-11.5,25,-11.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-11,21,-11</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-22.5,23,-11.5</points>
<intersection>-22.5 4</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23,-22.5,59.5,-22.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>23 3</intersection>
<intersection>34 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>34,-45.5,34,-22.5</points>
<intersection>-45.5 6</intersection>
<intersection>-22.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>34,-45.5,59.5,-45.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>34 5</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-8.5,45,-7.5</points>
<intersection>-8.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-8.5,59.5,-8.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection>
<intersection>53.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-7.5,45,-7.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53.5,-20.5,53.5,-8.5</points>
<intersection>-20.5 4</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53.5,-20.5,59.5,-20.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>53.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-33.5,44,-10.5</points>
<intersection>-33.5 4</intersection>
<intersection>-11.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-10.5,59.5,-10.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-11.5,44,-11.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>44,-33.5,59.5,-33.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-18.5,37.5,-12.5</points>
<intersection>-18.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-12.5,59.5,-12.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-18.5,37.5,-18.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-28,37.5,-24.5</points>
<intersection>-28 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-24.5,59.5,-24.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-28,37.5,-28</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-36,37,-35.5</points>
<intersection>-36 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-35.5,59.5,-35.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-36,37,-36</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-47.5,37,-47</points>
<intersection>-47.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-47.5,59.5,-47.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-47,37,-47</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-24,82,-10.5</points>
<intersection>-24 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-24,85.5,-24</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-10.5,82,-10.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-26,75.5,-22.5</points>
<intersection>-26 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-26,85.5,-26</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-22.5,75.5,-22.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-33.5,76,-28</points>
<intersection>-33.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-28,85.5,-28</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-33.5,76,-33.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-45.5,75.5,-36.5</points>
<intersection>-45.5 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-36.5,82.5,-36.5</points>
<intersection>75.5 0</intersection>
<intersection>82.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-45.5,75.5,-45.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-36.5,82.5,-30</points>
<intersection>-36.5 1</intersection>
<intersection>-30 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-30,85.5,-30</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>82.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-84.9016,37.4463,52.7984,-106.173</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>-38.5,24.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>-39,19.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>-35,-8</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-36.5,-19</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-38,-31</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-37,-41</position>
<gparam>LABEL_TEXT I4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>-37.5,13</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>-36.5,-54</position>
<gparam>LABEL_TEXT I5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-38,-66</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-37,-76</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>-38,-87</position>
<gparam>LABEL_TEXT I8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND4</type>
<position>66,-5.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND4</type>
<position>66,-17</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>31 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND4</type>
<position>66,-28</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>30 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND4</type>
<position>66,-39</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>29 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND4</type>
<position>66,-51</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>28 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND4</type>
<position>66,-62.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>27 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND4</type>
<position>66,-73.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>26 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND4</type>
<position>66,-84.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>25 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_OR4</type>
<position>92,-24.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>16 </input>
<input>
<ID>IN_3</ID>17 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR4</type>
<position>93,-74.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_OR2</type>
<position>123,-47</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>133.5,-47.5</position>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>-30.5,26.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>-30.5,22</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-30.5,13</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>-30,-8.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>-30,-20</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>-30.5,-31</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>-30.5,-42</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>-30,-54</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>-30,-65.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-30.5,-76.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>-30.5,-87.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_SMALL_INVERTER</type>
<position>-12,26.5</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_SMALL_INVERTER</type>
<position>-12,22</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_SMALL_INVERTER</type>
<position>-11,13</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-21.5,83,-5.5</points>
<intersection>-21.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-21.5,89,-21.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-5.5,83,-5.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-23.5,79,-17</points>
<intersection>-23.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-23.5,89,-23.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-17,79,-17</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-26.5,79,-25.5</points>
<intersection>-26.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-25.5,89,-25.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-26.5,79,-26.5</points>
<intersection>69 3</intersection>
<intersection>79 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-28,69,-26.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>-26.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-39,79,-27.5</points>
<intersection>-39 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-27.5,89,-27.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-39,79,-39</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-71.5,85,-51</points>
<intersection>-71.5 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-71.5,90,-71.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-51,85,-51</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-73.5,81,-62.5</points>
<intersection>-73.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-73.5,90,-73.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-62.5,81,-62.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-75.5,79.5,-73.5</points>
<intersection>-75.5 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-75.5,90,-75.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-73.5,79.5,-73.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-84.5,79.5,-77.5</points>
<intersection>-84.5 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-77.5,90,-77.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-84.5,79.5,-84.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-46,108,-24.5</points>
<intersection>-46 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-46,120,-46</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-24.5,108,-24.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-74.5,108.5,-48</points>
<intersection>-74.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-48,120,-48</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-74.5,108.5,-74.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-47.5,130,-47</points>
<intersection>-47.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-47.5,134.5,-47.5</points>
<connection>
<GID>66</GID>
<name>N_in1</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126,-47,130,-47</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,-87.5,63,-87.5</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,-76.5,63,-76.5</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-65.5,63,-65.5</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-54,63,-54</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,-42,63,-42</points>
<connection>
<GID>48</GID>
<name>IN_3</name></connection>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,-31,63,-31</points>
<connection>
<GID>46</GID>
<name>IN_3</name></connection>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-20,63,-20</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-8.5,63,-8.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,13,-13,13</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-14 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14,-85.5,-14,13</points>
<intersection>-85.5 10</intersection>
<intersection>-63.5 8</intersection>
<intersection>-40 6</intersection>
<intersection>-18 4</intersection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-14,-18,63,-18</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>-14 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-14,-40,63,-40</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>-14 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-14,-63.5,63,-63.5</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>-14 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-14,-85.5,63,-85.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>-14 3</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,22,-14,22</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19,-83.5,-19,22</points>
<intersection>-83.5 10</intersection>
<intersection>-61.5 8</intersection>
<intersection>-50 6</intersection>
<intersection>-27 4</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-19,-27,63,-27</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-19,-50,63,-50</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-19,-61.5,63,-61.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-19,-83.5,63,-83.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,26.5,-14,26.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-25.5,-81.5,-25.5,26.5</points>
<intersection>-81.5 5</intersection>
<intersection>-70.5 9</intersection>
<intersection>-59.5 11</intersection>
<intersection>-48 8</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-25.5,-81.5,63,-81.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-25.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-25.5,-48,63,-48</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-25.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-25.5,-70.5,63,-70.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-25.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-25.5,-59.5,63,-59.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-25.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-2.5,49,26.5</points>
<intersection>-2.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-2.5,63,-2.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,26.5,49,26.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-36,56,-2.5</points>
<intersection>-36 6</intersection>
<intersection>-25 7</intersection>
<intersection>-14 4</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-14,63,-14</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>56,-36,63,-36</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>56,-25,63,-25</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-4.5,26.5,22</points>
<intersection>-4.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-4.5,63,-4.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection>
<intersection>51.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,22,26.5,22</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51.5,-72.5,51.5,-4.5</points>
<intersection>-72.5 8</intersection>
<intersection>-38 6</intersection>
<intersection>-16 4</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51.5,-16,63,-16</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>51.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51.5,-38,63,-38</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>51.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>51.5,-72.5,63,-72.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>51.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-6.5,63,-6.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>7 3</intersection>
<intersection>46 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7,-6.5,7,13</points>
<intersection>-6.5 1</intersection>
<intersection>13 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-9,13,7,13</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>7 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>46,-74.5,46,-6.5</points>
<intersection>-74.5 10</intersection>
<intersection>-52 8</intersection>
<intersection>-29 6</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>46,-29,63,-29</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>46 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>46,-52,63,-52</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>46 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>46,-74.5,63,-74.5</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>46 5</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 2>
<page 3>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 3>
<page 4>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 4>
<page 5>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5308,122.4,-94.1308</PageViewport></page 9></circuit>