<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-17.1889,17.8889,61.3889,-64.0667</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>24,-5.5</position>
<gparam>LABEL_TEXT 2 to 4 line Decoder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>-9.5,-25</position>
<gparam>LABEL_TEXT A.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>31.5,-23.5</position>
<gparam>LABEL_TEXT D.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>-7,-14.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>39,-40</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>35,-33.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>39,-49</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-8,-18</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-8.5,-22.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>20,-24</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,-21.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>3,-26.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>27.5,-24</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>29.5,-34</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>22,-34</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>26,-40.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>34.5,-40.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>27.5,-49.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>34,-49.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-21.5,0,-18</points>
<intersection>-21.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-18,0,-18</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-21.5,2,-21.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-1.5 3</intersection>
<intersection>0 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-39.5,-1.5,-21.5</points>
<intersection>-39.5 4</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1.5,-39.5,23,-39.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-1.5 3</intersection>
<intersection>21.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>21.5,-48.5,21.5,-39.5</points>
<intersection>-48.5 6</intersection>
<intersection>-39.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-48.5,24.5,-48.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>21.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-23,11.5,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-23,17,-23</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-21.5,11.5,-21.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-33,17,-23</points>
<intersection>-33 4</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-33,19,-33</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>17 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-26.5,-3,-22.5</points>
<intersection>-26.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-22.5,-3,-22.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-3,-26.5,1,-26.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-3 0</intersection>
<intersection>-0.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-0.5,-35,-0.5,-26.5</points>
<intersection>-35 4</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-0.5,-35,24.5,-35</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-0.5 3</intersection>
<intersection>24.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>24.5,-50.5,24.5,-35</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-35 4</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-26.5,11,-25</points>
<intersection>-26.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-25,17,-25</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-1.5 3</intersection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-26.5,11,-26.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-41.5,-1.5,-25</points>
<intersection>-41.5 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1.5,-41.5,23,-41.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-1.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-24,26.5,-24</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-34,28.5,-34</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-40.5,33.5,-40.5</points>
<connection>
<GID>17</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-49.5,33,-49.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-17.1889,17.8889,61.3889,-64.0667</PageViewport>
<gate>
<ID>20</ID>
<type>AA_AND3</type>
<position>25.5,-19.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND3</type>
<position>25.5,-9</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND3</type>
<position>26,-30</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>22 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND3</type>
<position>26,-41</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND3</type>
<position>25.5,-49.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND3</type>
<position>26,-59</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND3</type>
<position>25.5,-69</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>22 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND3</type>
<position>25.5,-79</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>33,-9</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>33,-20</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>32,-30</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>32,-41</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>32,-49.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>32,-59</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>31.5,-69.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>32,-78.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>39,-8.5</position>
<gparam>LABEL_TEXT D.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>38.5,-19.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>39,-30</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>37.5,-40.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>38.5,-49</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>39,-58.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>39,-69.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>38.5,-78</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AE_SMALL_INVERTER</type>
<position>3.5,-9.5</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_SMALL_INVERTER</type>
<position>3.5,-5.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,0</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>-6.5,3</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>-8,-2.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-8,-8</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>-6.5,6.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>-12.5,-1</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>-9,-10.5</position>
<gparam>LABEL_TEXT A.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>24,13</position>
<gparam>LABEL_TEXT 3 to 8 line Decoder </gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-9,32,-9</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-20,30,-19.5</points>
<intersection>-20 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-19.5,30,-19.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-20,32,-20</points>
<connection>
<GID>29</GID>
<name>N_in0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-30,31,-30</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-41,31,-41</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<connection>
<GID>23</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-49.5,31,-49.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-59,31,-59</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>25</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-69,30.5,-69</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-69.5,30.5,-69</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-79,29.5,-78.5</points>
<intersection>-79 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-79,29.5,-79</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-78.5,31,-78.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,2,-3.5,3</points>
<intersection>2 2</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,3,-3.5,3</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-3.5,2,22.5,2</points>
<intersection>-3.5 0</intersection>
<intersection>2 5</intersection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-77,22.5,2</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-57 6</intersection>
<intersection>2 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>2,0,2,2</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22.5,-57,23,-57</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-5.5,-2.5,-2.5</points>
<intersection>-5.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-5.5,1.5,-5.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-2.5 0</intersection>
<intersection>-2 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-2.5,-2.5,-2.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2,-30,-2,-5.5</points>
<intersection>-30 4</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-2,-30,23,-30</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-2 3</intersection>
<intersection>23 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23,-69,23,-30</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-69 6</intersection>
<intersection>-30 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22.5,-69,23,-69</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>22.5 7</intersection>
<intersection>23 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>22.5,-79,22.5,-69</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-69 6</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-9.5,-2.5,-8</points>
<intersection>-9.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-9.5,1.5,-9.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-2.5 0</intersection>
<intersection>-1 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-8,-2.5,-8</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1,-21.5,-1,-9.5</points>
<intersection>-21.5 4</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1,-21.5,23,-21.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-1 3</intersection>
<intersection>23 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23,-81,23,-21.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<intersection>-81 7</intersection>
<intersection>-21.5 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-81,23,-81</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>23 5</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-7,14,0</points>
<intersection>-7 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,0,14,0</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-7,22.5,-7</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-28,22.5,-7</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-28 4</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-28,23,-28</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>22.5 3</intersection>
<intersection>23 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23,-39,23,-28</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-28 4</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-9,14,-5.5</points>
<intersection>-9 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-5.5,14,-5.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-9,22.5,-9</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-59,22.5,-9</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-59 6</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22.5,-59,23,-59</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-11,14,-9.5</points>
<intersection>-11 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-9.5,14,-9.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-11,23,-11</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>14 0</intersection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-51.5,23,-11</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-51.5 4</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-51.5,23,-51.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>22.5 5</intersection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>22.5,-71,22.5,-51.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>-51.5 4</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>