<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,44.2,-46.1</PageViewport>
<gate>
<ID>1</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-33</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>4,-24.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>11.5,-29.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>36,-26.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>35.5,-34</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>17,-13</position>
<gparam>LABEL_TEXT D  FLIP FLOP</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>BE_JKFF_LOW</type>
<position>24,-28.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>3 </output>
<input>
<ID>clock</ID>5 </input>
<output>
<ID>nQ</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>3.5,-21</position>
<gparam>LABEL_TEXT d</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>34,-23</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>12,-26.5</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>34.5,-30.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-33,6,-24.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-33 3</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-26.5,21,-26.5</points>
<connection>
<GID>7</GID>
<name>J</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6,-33,9.5,-33</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-33,17,-30.5</points>
<intersection>-33 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-33,17,-33</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-30.5,21,-30.5</points>
<connection>
<GID>7</GID>
<name>K</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-26.5,35,-26.5</points>
<connection>
<GID>7</GID>
<name>Q</name></connection>
<connection>
<GID>4</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-34,30.5,-30.5</points>
<intersection>-34 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-30.5,30.5,-30.5</points>
<connection>
<GID>7</GID>
<name>nQ</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-34,34.5,-34</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-29.5,21,-29.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>21 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>21,-29.5,21,-28.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>