<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,44.2,-46.1</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>5.5,-23</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>12,-35</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>9.5,-27</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>41.5,-27</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>41,-35.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>21.5,-11</position>
<gparam>LABEL_TEXT JK FLIP FLOP</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>6,-19.5</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>12.5,-24.5</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>13.5,-32</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>40.5,-23.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>40,-32</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>BE_JKFF_LOW</type>
<position>28.5,-26.5</position>
<input>
<ID>J</ID>4 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>2 </output>
<input>
<ID>clear</ID>1 </input>
<input>
<ID>clock</ID>1 </input>
<output>
<ID>nQ</ID>3 </output>
<input>
<ID>set</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-27,18.5,-26.5</points>
<intersection>-27 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-26.5,25.5,-26.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>18.5 0</intersection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-27,18.5,-27</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-30.5,23,-22.5</points>
<intersection>-30.5 5</intersection>
<intersection>-26.5 1</intersection>
<intersection>-22.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23,-30.5,28.5,-30.5</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>23 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>23,-22.5,28.5,-22.5</points>
<connection>
<GID>12</GID>
<name>set</name></connection>
<intersection>23 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-27,36,-24.5</points>
<intersection>-27 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-27,40.5,-27</points>
<connection>
<GID>4</GID>
<name>N_in0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-24.5,36,-24.5</points>
<connection>
<GID>12</GID>
<name>Q</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-35.5,35,-28.5</points>
<intersection>-35.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-28.5,35,-28.5</points>
<connection>
<GID>12</GID>
<name>nQ</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-35.5,40,-35.5</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-24.5,16.5,-23</points>
<intersection>-24.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-23,16.5,-23</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-24.5,25.5,-24.5</points>
<connection>
<GID>12</GID>
<name>J</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-35,19.5,-28.5</points>
<intersection>-35 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-28.5,25.5,-28.5</points>
<connection>
<GID>12</GID>
<name>K</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-35,19.5,-35</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>