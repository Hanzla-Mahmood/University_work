<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-20.4788,-0.178221,122.517,-75.5316</PageViewport>
<gate>
<ID>2</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-15</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>6.5,-5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_SMALL_INVERTER</type>
<position>16,-21.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>16.5,-29.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>6.5,-12.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>6.5,-9</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>6.5,-16</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>6,-20</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>7,-24</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>7.5,-31</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>8.5,-34</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>74.5,-13</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR4</type>
<position>42,-17.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>10 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>80.5,-13</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>30,-20</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>28.5,-29</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>81,-28</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>75,-28.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR3</type>
<position>43.5,-34</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>62.5,-49</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>27,-38</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>26.5,-44</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>76,-59.5</position>
<gparam>LABEL_TEXT d</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AE_OR3</type>
<position>44.5,-49.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>1 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>58.5,-49.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>58.5,-84</position>
<gparam>LABEL_TEXT e</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AE_OR3</type>
<position>45,-59.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>74.5,-96.5</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AE_OR3</type>
<position>57.5,-59.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>23 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>79,-116.5</position>
<gparam>LABEL_TEXT g</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>71,-59.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>33,-58</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>33.5,-64.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>44,-66.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND3</type>
<position>39,-74</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>1 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_OR2</type>
<position>46,-84</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>31,-83.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>31.5,-90</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>54,-84</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>75,-117</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>71,-96.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR4</type>
<position>37,-101</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>23.5,-97.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>22.5,-104</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>23.5,-111.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_OR4</type>
<position>31.5,-136</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<input>
<ID>IN_2</ID>34 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>10,-133</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>11,-139.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>-1,-143</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-32,14.5,-29.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-32,25.5,-32</points>
<intersection>14.5 0</intersection>
<intersection>24 6</intersection>
<intersection>25.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-31,14.5,-31</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25.5,-32,25.5,-30</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>24,-51.5,24,-32</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-51.5 7</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>24,-51.5,41.5,-51.5</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>24 6</intersection>
<intersection>36 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>36,-76,36,-51.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>-51.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-17.5,65,-13</points>
<intersection>-17.5 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-13,73.5,-13</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-17.5,65,-17.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-14.5,23.5,-9</points>
<intersection>-14.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-9,23.5,-9</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-14.5,42,-14.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection>
<intersection>42 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42,-104,42,-14.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-104 4</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28.5,-104,42,-104</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>28.5 5</intersection>
<intersection>42 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>28.5,-139,28.5,-104</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>-138.5 6</intersection>
<intersection>-104 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>8,-138.5,28.5,-138.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>28.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-20,35,-18.5</points>
<intersection>-20 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-18.5,39,-18.5</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-20,35,-20</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-40.5,34,-16.5</points>
<intersection>-40.5 4</intersection>
<intersection>-24 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-24,34,-24</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>13.5 3</intersection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-16.5,39,-16.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-24,13.5,-21.5</points>
<intersection>-24 1</intersection>
<intersection>-21.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-40.5,34,-40.5</points>
<intersection>24 5</intersection>
<intersection>30 7</intersection>
<intersection>34 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>24,-40.5,24,-39</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13.5,-21.5,14,-21.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>30,-89,30,-40.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-89 9</intersection>
<intersection>-63.5 8</intersection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>30,-63.5,30.5,-63.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>30 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>8,-89,30,-89</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>8 10</intersection>
<intersection>30 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>8,-142,8,-89</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-142 11</intersection>
<intersection>-89 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-4,-142,8,-142</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>8 10</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-19,24,-15</points>
<intersection>-19 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-15,24,-15</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-19,27,-19</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-32,24.5,-19</points>
<intersection>-32 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-32,40.5,-32</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection>
<intersection>30.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30.5,-82.5,30.5,-32</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>-82.5 7</intersection>
<intersection>-65.5 6</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30.5,-65.5,41,-65.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>30.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>28,-82.5,30.5,-82.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>30.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-21</points>
<intersection>-29.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-29.5,24,-29.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>23.5 3</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-21,27,-21</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-59,23.5,-29.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-59 4</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23.5,-59,30,-59</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>23.5 3</intersection>
<intersection>24.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>24.5,-67.5,24.5,-59</points>
<intersection>-67.5 7</intersection>
<intersection>-59 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>24.5,-67.5,41,-67.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>24.5 6</intersection>
<intersection>28 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>28,-98.5,28,-67.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-98.5 10</intersection>
<intersection>-91 9</intersection>
<intersection>-67.5 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>28,-91,28.5,-91</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>28 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>20.5,-98.5,28,-98.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>20.5 11</intersection>
<intersection>28 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>20.5,-144,20.5,-98.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-144 12</intersection>
<intersection>-98.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-4,-144,20.5,-144</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>20.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-29,35,-20.5</points>
<intersection>-29 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-20.5,39,-20.5</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-29,35,-29</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-34,60,-28.5</points>
<intersection>-34 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-28.5,74,-28.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-34,60,-34</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-28,17,-15</points>
<intersection>-28 2</intersection>
<intersection>-16 1</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-16,17,-16</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-28,41.5,-28</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection>
<intersection>41.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>17,-15,18.5,-15</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>41.5,-72,41.5,-28</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-72 5</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>19.5,-72,41.5,-72</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>19.5 6</intersection>
<intersection>41.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>19.5,-134,19.5,-72</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-134 8</intersection>
<intersection>-110.5 7</intersection>
<intersection>-72 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>19.5,-110.5,20.5,-110.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>19.5 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-134,19.5,-134</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>19.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-38,35,-34</points>
<intersection>-38 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-38,35,-38</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-34,40.5,-34</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-44,35,-36</points>
<intersection>-44 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-36,40.5,-36</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-44,35,-44</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-49.5,20.5,-22</points>
<intersection>-49.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-22,20.5,-22</points>
<intersection>18 3</intersection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-49.5,41.5,-49.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection>
<intersection>23.5 5</intersection>
<intersection>36 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-22,18,-21.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>23.5,-49.5,23.5,-45</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>36,-96.5,36,-49.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-96.5 7</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>19.5,-96.5,36,-96.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>19.5 8</intersection>
<intersection>36 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>19.5,-132,19.5,-96.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-132 9</intersection>
<intersection>-96.5 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>7,-132,19.5,-132</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>19.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-49.5,57.5,-49.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-59.5,70,-59.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-59.5,39,-58</points>
<intersection>-59.5 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-59.5,42,-59.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-58,39,-58</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-64.5,39,-61.5</points>
<intersection>-64.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-64.5,39,-64.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-61.5,42,-61.5</points>
<connection>
<GID>36</GID>
<name>IN_2</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-59.5,51,-57.5</points>
<intersection>-59.5 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-59.5,51,-59.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-57.5,54.5,-57.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-66.5,50.5,-59.5</points>
<intersection>-66.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-59.5,54.5,-59.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-66.5,50.5,-66.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-74,48,-61.5</points>
<intersection>-74 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-61.5,54.5,-61.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-74,48,-74</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-83.5,38.5,-83</points>
<intersection>-83.5 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-83,43,-83</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-83.5,38.5,-83.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-90,38.5,-85</points>
<intersection>-90 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-85,43,-85</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-90,38.5,-90</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-84,53,-84</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-101,55.5,-96.5</points>
<intersection>-101 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-96.5,70,-96.5</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-101,55.5,-101</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-98,30.5,-97.5</points>
<intersection>-98 1</intersection>
<intersection>-97.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-98,34,-98</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-97.5,30.5,-97.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-104,29.5,-100</points>
<intersection>-104 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-100,34,-100</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-104,29.5,-104</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-111.5,30,-102</points>
<intersection>-111.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-102,34,-102</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-111.5,30,-111.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-136,54.5,-117</points>
<intersection>-136 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-117,74,-117</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-136,54.5,-136</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-133,28.5,-133</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-139.5,21,-135</points>
<intersection>-139.5 2</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-135,28.5,-135</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-139.5,21,-139.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-143,15,-137</points>
<intersection>-143 2</intersection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-137,28.5,-137</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-143,15,-143</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 1>
<page 2>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 2>
<page 3>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 3>
<page 4>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 4>
<page 5>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 5>
<page 6>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 6>
<page 7>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 7>
<page 8>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 8>
<page 9>
<PageViewport>0,31.5808,338.954,-147.035</PageViewport></page 9></circuit>