<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-53.4083,-12.1568,164.192,-119.712</PageViewport>
<gate>
<ID>2</ID>
<type>AE_OR4</type>
<position>71.5,-64</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND4</type>
<position>44,-48</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND4</type>
<position>44,-62.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND4</type>
<position>44.5,-73</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>7 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND4</type>
<position>44,-83.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>9,-51</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>8.5,-65.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>8.5,-76</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>10.5,-86.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>0.5,-27.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>0,-34.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>0,-41</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_SMALL_INVERTER</type>
<position>6,-27.5</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,-34.5</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_SMALL_INVERTER</type>
<position>6.5,-41</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>76.5,-64</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-3.5,-26.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-3,-33.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>-3.5,-40.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>10,-54</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>9.5,-68</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>9.5,-78</position>
<gparam>LABEL_TEXT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>10.5,-88.5</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-61,57.5,-48</points>
<intersection>-61 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-48,57.5,-48</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-61,68.5,-61</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-63,57.5,-62.5</points>
<intersection>-63 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-62.5,57.5,-62.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-63,68.5,-63</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-73,58,-65</points>
<intersection>-73 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-73,58,-73</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58,-65,68.5,-65</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-83.5,57.5,-67</points>
<intersection>-83.5 1</intersection>
<intersection>-67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-83.5,57.5,-83.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-67,68.5,-67</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-51,41,-51</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-65.5,41,-65.5</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-76,41.5,-76</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-86.5,41,-86.5</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-64,75.5,-64</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>29</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-45,24.5,-27.5</points>
<intersection>-45 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-45,41,-45</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection>
<intersection>34 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-27.5,24.5,-27.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-59.5,34,-45</points>
<intersection>-59.5 4</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34,-59.5,41,-59.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-47,25,-34.5</points>
<intersection>-47 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-47,41,-47</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection>
<intersection>26.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-34.5,25,-34.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-72,26.5,-47</points>
<intersection>-72 4</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-72,41.5,-72</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-27.5,33,-27.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-70,33,-27.5</points>
<intersection>-70 4</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-70,41.5,-70</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection>
<intersection>35.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35.5,-80.5,35.5,-70</points>
<intersection>-80.5 6</intersection>
<intersection>-70 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-80.5,41,-80.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>35.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-34.5,5.5,-34.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>4.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-61.5,4.5,-34.5</points>
<intersection>-61.5 4</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>4.5,-61.5,41,-61.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>4.5 3</intersection>
<intersection>41 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>41,-82.5,41,-61.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-61.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-41,4.5,-41</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>3 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3,-63.5,3,-41</points>
<intersection>-63.5 5</intersection>
<intersection>-49 6</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>3,-63.5,41,-63.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>3 3</intersection>
<intersection>39 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>3,-49,41,-49</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>3 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>39,-74,39,-63.5</points>
<intersection>-74 8</intersection>
<intersection>-63.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>39,-74,41.5,-74</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>39 7</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-84.5,24.5,-41</points>
<intersection>-84.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-41,24.5,-41</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-84.5,41,-84.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>