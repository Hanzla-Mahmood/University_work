<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-17.1889,17.8889,61.3889,-64.0667</PageViewport>
<gate>
<ID>1</ID>
<type>BE_JKFF_LOW_NT</type>
<position>12,-29.5</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>3 </input>
<output>
<ID>Q</ID>4 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>24,-29.5</position>
<input>
<ID>J</ID>4 </input>
<input>
<ID>K</ID>4 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>BE_JKFF_LOW_NT</type>
<position>36.5,-30</position>
<input>
<ID>J</ID>6 </input>
<input>
<ID>K</ID>6 </input>
<output>
<ID>Q</ID>7 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>BB_CLOCK</type>
<position>0.5,-35.5</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-1,-17.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-20.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>25.5,-17</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>43,-24.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>18,-3.5</position>
<gparam>LABEL_TEXT 3-Bit Synchronous Counter</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-35.5,31,-35.5</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<intersection>6 5</intersection>
<intersection>18 4</intersection>
<intersection>31 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>18,-35.5,18,-29.5</points>
<intersection>-35.5 1</intersection>
<intersection>-29.5 9</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>6,-35.5,6,-29.5</points>
<intersection>-35.5 1</intersection>
<intersection>-29.5 10</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>31,-35.5,31,-30</points>
<intersection>-35.5 1</intersection>
<intersection>-30 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>31,-30,33.5,-30</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>31 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>18,-29.5,21,-29.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>18 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>6,-29.5,9,-29.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>6 5</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-27.5,5,-17.5</points>
<intersection>-27.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-27.5,9,-27.5</points>
<connection>
<GID>1</GID>
<name>J</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-17.5,5,-17.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-31.5,3,-20.5</points>
<intersection>-31.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-31.5,9,-31.5</points>
<connection>
<GID>1</GID>
<name>K</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-20.5,3,-20.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-27.5,21,-27.5</points>
<connection>
<GID>2</GID>
<name>J</name></connection>
<connection>
<GID>1</GID>
<name>Q</name></connection>
<intersection>18 5</intersection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-31.5,20,-27.5</points>
<intersection>-31.5 4</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-31.5,21,-31.5</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>18,-27.5,18,-16</points>
<intersection>-27.5 1</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>18,-16,22.5,-16</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>18 5</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-27.5,27,-21</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,-21,27,-21</points>
<intersection>22 3</intersection>
<intersection>27 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-21,22,-18</points>
<intersection>-21 2</intersection>
<intersection>-18 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22,-18,22.5,-18</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>22 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-28,30.5,-17</points>
<intersection>-28 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-28,33.5,-28</points>
<connection>
<GID>3</GID>
<name>J</name></connection>
<intersection>30.5 0</intersection>
<intersection>32 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-17,30.5,-17</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-32,32,-28</points>
<intersection>-32 4</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,-32,33.5,-32</points>
<connection>
<GID>3</GID>
<name>K</name></connection>
<intersection>32 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-28,40.5,-24.5</points>
<intersection>-28 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-24.5,42,-24.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-28,40.5,-28</points>
<connection>
<GID>3</GID>
<name>Q</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>