<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-15,18,107.4,-46.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>24.5,-16</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>23,-29.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BE_NOR2</type>
<position>51.5,-17</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BE_NOR2</type>
<position>51.5,-28.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>8.5,-15</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>5.5,-23</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>8,-30.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>60.5,-28.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>58.5,-17</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>7.5,-12</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>7,-26.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>5,-19</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>60.5,-13</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>62,-25.5</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>30,6</position>
<gparam>LABEL_TEXT SR Flip Flop using NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-16,48.5,-16</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-29.5,48.5,-29.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-28.5,20,-17</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-17,21.5,-17</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-23,20,-23</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-15,21.5,-15</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>21.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>21.5,-15,21.5,-15</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-30.5,20,-30.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>20 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>20,-30.5,20,-30.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-17,57.5,-17</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55.5,-23.5,55.5,-17</points>
<intersection>-23.5 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48.5,-23.5,55.5,-23.5</points>
<intersection>48.5 7</intersection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>48.5,-27.5,48.5,-23.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-23.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-28.5,46,-18</points>
<intersection>-28.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-28.5,59.5,-28.5</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-18,48.5,-18</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-64.5</PageViewport></page 9></circuit>