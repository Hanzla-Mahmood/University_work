<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>10.5413,-0.743451,70.8678,-63.6632</PageViewport>
<gate>
<ID>1</ID>
<type>AI_XOR2</type>
<position>31.5,-26</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>253,-48</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>49,-30</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>32.5,-37</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>63.5,-44.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>17.5,-25</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>18,-30</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>25.5,-41</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>60,-15.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>53.5,-34.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>14.5,-24.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>15,-29.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>23.5,-40</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>47.5,-26</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>52.5,-48</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>90.5,-27</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AI_XOR2</type>
<position>108,-31</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>91.5,-38</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>122.5,-45.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>76.5,-26</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>77,-31</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>119,-16.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>112.5,-35.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>73.5,-25.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>74,-30.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>106.5,-27</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>111.5,-49</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AI_XOR2</type>
<position>151.5,-28.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AI_XOR2</type>
<position>169,-32.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>152.5,-39.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>183.5,-47</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>137.5,-27.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>138,-32.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>180,-18</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>173.5,-37</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>134.5,-27</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>135,-32</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>167.5,-28.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>172.5,-50.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>210,-29.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AI_XOR2</type>
<position>227.5,-33.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>211,-40.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_OR2</type>
<position>242,-48</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>196,-28.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>196.5,-33.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>238.5,-19</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>232,-38</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>193,-28</position>
<gparam>LABEL_TEXT A4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>193,-33</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>226,-29.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>231,-51.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>38,-14.5</position>
<gparam>LABEL_TEXT Ripple Carry Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-25,28.5,-25</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-36,24,-25</points>
<intersection>-36 4</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-36,29.5,-36</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-38,23,-27</points>
<intersection>-38 3</intersection>
<intersection>-30 4</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-27,28.5,-27</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23,-38,29.5,-38</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>20,-30,23,-30</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245,-48,252,-48</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-30,56,-15.5</points>
<intersection>-30 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-15.5,59,-15.5</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-30,56,-30</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-33.5,40,-26</points>
<intersection>-33.5 3</intersection>
<intersection>-29 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-29,46,-29</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-26,40,-26</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40,-33.5,50.5,-33.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-41,36,-31</points>
<intersection>-41 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-31,46,-31</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection>
<intersection>42 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-41,36,-41</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42,-35.5,42,-31</points>
<intersection>-35.5 4</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42,-35.5,50.5,-35.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>42 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-45.5,40,-37</points>
<intersection>-45.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-45.5,60.5,-45.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-37,40,-37</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-43.5,59,-34.5</points>
<intersection>-43.5 4</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-34.5,59,-34.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>59,-43.5,60.5,-43.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-26,87.5,-26</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>82.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-37,82.5,-26</points>
<intersection>-37 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-37,88.5,-37</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>82.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-39,82,-28</points>
<intersection>-39 3</intersection>
<intersection>-31 4</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-28,87.5,-28</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>82,-39,88.5,-39</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>79,-31,82,-31</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-31,115,-16.5</points>
<intersection>-31 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-16.5,118,-16.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-31,115,-31</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-34.5,99,-27</points>
<intersection>-34.5 3</intersection>
<intersection>-30 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-30,105,-30</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-27,99,-27</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99,-34.5,109.5,-34.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-32,105,-32</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>101 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101,-44.5,101,-32</points>
<intersection>-44.5 5</intersection>
<intersection>-36.5 4</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>101,-36.5,109.5,-36.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>101 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-44.5,101,-44.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>101 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-46.5,99,-38</points>
<intersection>-46.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-46.5,119.5,-46.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-38,99,-38</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-44.5,118,-35.5</points>
<intersection>-44.5 4</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-35.5,118,-35.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>118,-44.5,119.5,-44.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,-27.5,148.5,-27.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>144 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>144,-38.5,144,-27.5</points>
<intersection>-38.5 4</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>144,-38.5,149.5,-38.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>144 3</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-40.5,143,-29.5</points>
<intersection>-40.5 3</intersection>
<intersection>-32.5 4</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-29.5,148.5,-29.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>143,-40.5,149.5,-40.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>140,-32.5,143,-32.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-32.5,176,-18</points>
<intersection>-32.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-18,179,-18</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-32.5,176,-32.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-36,160,-28.5</points>
<intersection>-36 3</intersection>
<intersection>-31.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-31.5,166,-31.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154.5,-28.5,160,-28.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>160,-36,170.5,-36</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-33.5,166,-33.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>162 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>162,-45.5,162,-33.5</points>
<intersection>-45.5 5</intersection>
<intersection>-38 4</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>162,-38,170.5,-38</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>162 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>125.5,-45.5,162,-45.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>162 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-48,160,-39.5</points>
<intersection>-48 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-48,180.5,-48</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-39.5,160,-39.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-46,179,-37</points>
<intersection>-46 4</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>176.5,-37,179,-37</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>179,-46,180.5,-46</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-28.5,207,-28.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>203 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>203,-39.5,203,-28.5</points>
<intersection>-39.5 4</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>203,-39.5,208,-39.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>203 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-41.5,201.5,-30.5</points>
<intersection>-41.5 3</intersection>
<intersection>-33.5 4</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201.5,-30.5,207,-30.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>201.5,-41.5,208,-41.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198.5,-33.5,201.5,-33.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-33.5,234.5,-19</points>
<intersection>-33.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,-19,237.5,-19</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>230.5,-33.5,234.5,-33.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-37,218.5,-29.5</points>
<intersection>-37 3</intersection>
<intersection>-32.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-32.5,224.5,-32.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213,-29.5,218.5,-29.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>218.5,-37,229,-37</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,-34.5,224.5,-34.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>220.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>220.5,-47,220.5,-34.5</points>
<intersection>-47 5</intersection>
<intersection>-39 4</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>220.5,-39,229,-39</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>220.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>186.5,-47,220.5,-47</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>220.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-49,218.5,-40.5</points>
<intersection>-49 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-49,239,-49</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-40.5,218.5,-40.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-47,237.5,-38</points>
<intersection>-47 4</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>235,-38,237.5,-38</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>237.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>237.5,-47,239,-47</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 1>
<page 2>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 2>
<page 3>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 3>
<page 4>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 4>
<page 5>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 5>
<page 6>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 6>
<page 7>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 7>
<page 8>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 8>
<page 9>
<PageViewport>0,121.035,338.954,-232.489</PageViewport></page 9></circuit>