<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-7.36667,7.66667,51.5667,-53.8</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>24,-7</position>
<gparam>LABEL_TEXT 4 to 2 Encoder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>1,-19</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>1.5,-25.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>2,-31.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>-2.5,-31</position>
<gparam>LABEL_TEXT E1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-3.5,-24.5</position>
<gparam>LABEL_TEXT E2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-4.5,-17.5</position>
<gparam>LABEL_TEXT E3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>40,-25</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>22.5,-22.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>21.5,-36</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>35.5,-37</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>45.5,-25</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>42,-36.5</position>
<gparam>LABEL_TEXT A.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-21.5,10,-19</points>
<intersection>-21.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-21.5,19.5,-21.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection>
<intersection>18.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-19,10,-19</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18.5,-35,18.5,-21.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-25.5,10,-23.5</points>
<intersection>-25.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-25.5,10,-25.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-23.5,19.5,-23.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-25,32,-22.5</points>
<intersection>-25 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-25,39,-25</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-22.5,32,-22.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-37,11,-31.5</points>
<intersection>-37 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-31.5,11,-31.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-37,18.5,-37</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-37,29.5,-36</points>
<intersection>-37 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-36,29.5,-36</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-37,34.5,-37</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>