<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-33.9125,31.4324,288.587,-127.973</PageViewport>
<gate>
<ID>1</ID>
<type>AI_XOR2</type>
<position>25.5,-17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>247,-39.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>43,-21.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>26.5,-28.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>57.5,-36</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>11.5,-16.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>12,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>19.5,-32.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>54,-7</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>47.5,-26</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>8.5,-16</position>
<gparam>LABEL_TEXT a1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>9,-21</position>
<gparam>LABEL_TEXT b1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>17.5,-31.5</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>41.5,-17.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>46.5,-39.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>84.5,-18.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AI_XOR2</type>
<position>102,-22.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>85.5,-29.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>116.5,-37</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>70.5,-17.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>71,-22.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>113,-8</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>106.5,-27</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>67.5,-17</position>
<gparam>LABEL_TEXT a2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>68,-22</position>
<gparam>LABEL_TEXT b2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>100.5,-18.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>105.5,-40.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AI_XOR2</type>
<position>145.5,-20</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AI_XOR2</type>
<position>163,-24</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>146.5,-31</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>177.5,-38.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>131.5,-19</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>132,-24</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>174,-9.5</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>167.5,-28.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>128.5,-18.5</position>
<gparam>LABEL_TEXT a3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>129,-23.5</position>
<gparam>LABEL_TEXT b3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>161.5,-20</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>166.5,-42</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>204,-21</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AI_XOR2</type>
<position>221.5,-25</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>205,-32</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_OR2</type>
<position>236,-39.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>190,-20</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>190.5,-25</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>232.5,-10.5</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>226,-29.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>187,-19.5</position>
<gparam>LABEL_TEXT a4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>187.5,-24.5</position>
<gparam>LABEL_TEXT b4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>220,-21</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>225,-43</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>117.5,-61.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_OR2</type>
<position>124.5,-88.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND2</type>
<position>178.5,-56</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_OR2</type>
<position>186,-80.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>123.5,-38</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>186,-39</position>
<input>
<ID>N_in2</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-16.5,22.5,-16.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-27.5,19,-16.5</points>
<intersection>-27.5 4</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-27.5,23.5,-27.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-29.5,17,-18.5</points>
<intersection>-29.5 3</intersection>
<intersection>-21.5 4</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-18.5,22.5,-18.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>17,-29.5,23.5,-29.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>14,-21.5,17,-21.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239,-39.5,246,-39.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-21.5,50,-7</points>
<intersection>-21.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-7,53,-7</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-21.5,50,-21.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-25,34,-17.5</points>
<intersection>-25 3</intersection>
<intersection>-20.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-20.5,40,-20.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-17.5,34,-17.5</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>34,-25,44.5,-25</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-32.5,30,-22.5</points>
<intersection>-32.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-22.5,40,-22.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection>
<intersection>36 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-32.5,30,-32.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-27,36,-22.5</points>
<intersection>-27 4</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-27,44.5,-27</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-37,34,-28.5</points>
<intersection>-37 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-37,54.5,-37</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-28.5,34,-28.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-35,53,-26</points>
<intersection>-35 4</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-26,53,-26</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53,-35,54.5,-35</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-17.5,81.5,-17.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-28.5,77.5,-17.5</points>
<intersection>-28.5 4</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>77.5,-28.5,82.5,-28.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-30.5,76,-19.5</points>
<intersection>-30.5 3</intersection>
<intersection>-22.5 4</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-19.5,81.5,-19.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>76,-30.5,82.5,-30.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73,-22.5,76,-22.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-22.5,109,-8</points>
<intersection>-22.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-8,112,-8</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-22.5,109,-22.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-26,93,-18.5</points>
<intersection>-26 3</intersection>
<intersection>-21.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-21.5,99,-21.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-18.5,93,-18.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>91,-26,103.5,-26</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>91 4</intersection>
<intersection>93 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91,-60.5,91,-26</points>
<intersection>-60.5 5</intersection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91,-60.5,114.5,-60.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>91 4</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-23.5,99,-23.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-62.5,84.5,-23.5</points>
<intersection>-62.5 6</intersection>
<intersection>-36 5</intersection>
<intersection>-28 4</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>84.5,-28,103.5,-28</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>84.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>60.5,-36,84.5,-36</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>84.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-62.5,114.5,-62.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>84.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-89.5,93,-29.5</points>
<intersection>-89.5 4</intersection>
<intersection>-38 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-38,113.5,-38</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-29.5,93,-29.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>93,-89.5,121.5,-89.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-36,112,-27</points>
<intersection>-36 4</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-27,112,-27</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112,-36,113.5,-36</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-19,142.5,-19</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>139 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>139,-30,139,-19</points>
<intersection>-30 4</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>139,-30,143.5,-30</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>139 3</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-32,137,-21</points>
<intersection>-32 3</intersection>
<intersection>-24 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-21,142.5,-21</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>137,-32,143.5,-32</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>134,-24,137,-24</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-24,170,-9.5</points>
<intersection>-24 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-9.5,173,-9.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-24,170,-24</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-27.5,154,-20</points>
<intersection>-27.5 3</intersection>
<intersection>-23 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-23,160,-23</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-20,154,-20</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>154,-27.5,164.5,-27.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection>
<intersection>157.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>157.5,-55,157.5,-27.5</points>
<intersection>-55 5</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>157.5,-55,175.5,-55</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>157.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-81.5,154,-31</points>
<intersection>-81.5 4</intersection>
<intersection>-39.5 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-39.5,174.5,-39.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149.5,-31,154,-31</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>154,-81.5,183,-81.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-37.5,173,-28.5</points>
<intersection>-37.5 4</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-28.5,173,-28.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>173,-37.5,174.5,-37.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192,-20,201,-20</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>198 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>198,-31,198,-20</points>
<intersection>-31 4</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>198,-31,202,-31</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>198 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-33,195.5,-22</points>
<intersection>-33 3</intersection>
<intersection>-25 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,-22,201,-22</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>195.5,-33,202,-33</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>192.5,-25,195.5,-25</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-25,228.5,-10.5</points>
<intersection>-25 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,-10.5,231.5,-10.5</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>224.5,-25,228.5,-25</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,-28.5,212.5,-21</points>
<intersection>-28.5 3</intersection>
<intersection>-24 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-24,218.5,-24</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-21,212.5,-21</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>212.5,-28.5,223,-28.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>212.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,-40.5,212.5,-32</points>
<intersection>-40.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212.5,-40.5,233,-40.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208,-32,212.5,-32</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>212.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-38.5,231.5,-29.5</points>
<intersection>-38.5 4</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>229,-29.5,231.5,-29.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>231.5,-38.5,233,-38.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-87.5,120.5,-61.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-87.5,121.5,-87.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-88.5,149.5,-29.5</points>
<intersection>-88.5 2</intersection>
<intersection>-57 4</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-29.5,164.5,-29.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection>
<intersection>160 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-88.5,149.5,-88.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>149.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>160,-29.5,160,-25</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>149.5,-57,175.5,-57</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-79.5,182,-56</points>
<intersection>-79.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-56,182,-56</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182,-79.5,183,-79.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-80.5,203.5,-26</points>
<intersection>-80.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203.5,-26,218.5,-26</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>203.5 0</intersection>
<intersection>215 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-80.5,203.5,-80.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>215,-30.5,215,-26</points>
<intersection>-30.5 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>215,-30.5,223,-30.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>215 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-38,121,-37</points>
<intersection>-38 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-38,122.5,-38</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-37,121,-37</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-40,186,-38.5</points>
<connection>
<GID>63</GID>
<name>N_in2</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,-38.5,186,-38.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>